module tb();
reg clk,rst;
wire Jrsel,sel31,selPc,regwrite,RegDst,MemRead,MemWrite,MemToReg,zero,PCsel,ALUSrcA,IRWrite,IorD;
wire [2:0] ALU_operation;
wire [1:0] alu_op,PCSrc,ALUSrcB;
wire [5:0] OPC,Func;
mips MIPS(clk,rst,Jrsel,sel31,selPc,ALU_operation,PCsel,ALUSrcA,ALUSrcB,RegDst,MemToReg,IRWrite,MemRead,MemWrite,IorD,regwrite,PCSrc,zero,OPC,Func);
controller CONTROLLER(clk,rst,zero,selPc,OPC,sel31,regwrite,RegDst,alu_op,MemRead,MemWrite,MemToReg,IorD,IRWrite,ALUSrcA,ALUSrcB,PCSrc,PCsel,Jrsel);
ALU_controller ALU_CONTROLLER(clk,alu_op,Func,ALU_operation);

initial begin
    #10 rst = 1;
    #20 rst = 0; 
    #20 clk=0;  
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;
    #20 clk=1;
    #20 clk=0;


end
endmodule